interface iface(input bit clk, rst);
  
  bit data_in;
  bit full;
 
endinterface: iface